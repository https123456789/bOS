<svg version="1.1" width="100%" height="100%" xmlns="http://www.w3.org/2000/svg">
	<defs>
		<radialGradient id="grad1" x1="0%" y1="0%" x2="100%" y2="0%">
			<stop offset="0%" style="stop-color: rgb(255, 255, 255);"></stop>
			<stop offset="100%" stlye="stop-color: rgb(0, 0, 0);"></stop>
		</radialGradient>
	</defs>
	<rect width="100%" height="100%" fill="url(#grad1)"></rect>
</svg>